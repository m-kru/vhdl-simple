library ieee;
   use ieee.std_logic_1164.all;

package simple is

   type t_slv_vector is array(natural range <>) of std_logic_vector;

end package;
